// array.pl 25 25 
// $Id: array.pl,v 1.5 2015-04-03 09:31:09 a Exp $ 
// Date: Sat Jul 11 17:31:06 2015
// AUTHOR: (C) moshahmed/at/gmail

module u(clock,enable,reset,set,in1,in2,out1,out2);
    input  clock,enable,reset,set,in1,in2;
    output out1,out2;
    reg    out1,out2;
    always@(posedge clock) begin
        if( enable )
            out1 <=in1;
        if( reset )
            out2 <= 0;
        else if( set )
            out2 <= 1;
        else if( enable )
            out2 <=in2;
        end
endmodule

module array(clock,enable,reset,set,
  in_00_01, ou_00_00, in_00_02, ou_00_01, in_00_03, ou_00_02, in_00_04, ou_00_03,  
  in_00_05, ou_00_04, in_00_06, ou_00_05, in_00_07, ou_00_06, in_00_08, ou_00_07,  
  in_00_09, ou_00_08, in_00_10, ou_00_09, in_00_11, ou_00_10, in_00_12, ou_00_11,  
  in_00_13, ou_00_12, in_00_14, ou_00_13, in_00_15, ou_00_14, in_00_16, ou_00_15,  
  in_00_17, ou_00_16, in_00_18, ou_00_17, in_00_19, ou_00_18, in_00_20, ou_00_19,  
  in_00_21, ou_00_20, in_00_22, ou_00_21, in_00_23, ou_00_22, in_00_24, ou_00_23,  
  in_00_25, ou_00_24, in_25_01, ou_25_01, in_25_02, ou_25_02, in_25_03, ou_25_03,  
  in_25_04, ou_25_04, in_25_05, ou_25_05, in_25_06, ou_25_06, in_25_07, ou_25_07,  
  in_25_08, ou_25_08, in_25_09, ou_25_09, in_25_10, ou_25_10, in_25_11, ou_25_11,  
  in_25_12, ou_25_12, in_25_13, ou_25_13, in_25_14, ou_25_14, in_25_15, ou_25_15,  
  in_25_16, ou_25_16, in_25_17, ou_25_17, in_25_18, ou_25_18, in_25_19, ou_25_19,  
  in_25_20, ou_25_20, in_25_21, ou_25_21, in_25_22, ou_25_22, in_25_23, ou_25_23,  
  in_25_24, ou_25_24, in_25_25, ou_25_25
);

input clock,enable,reset,set, 
  in_00_01, ou_00_00, in_00_02, ou_00_01, in_00_03, ou_00_02, in_00_04, ou_00_03,  
  in_00_05, ou_00_04, in_00_06, ou_00_05, in_00_07, ou_00_06, in_00_08, ou_00_07,  
  in_00_09, ou_00_08, in_00_10, ou_00_09, in_00_11, ou_00_10, in_00_12, ou_00_11,  
  in_00_13, ou_00_12, in_00_14, ou_00_13, in_00_15, ou_00_14, in_00_16, ou_00_15,  
  in_00_17, ou_00_16, in_00_18, ou_00_17, in_00_19, ou_00_18, in_00_20, ou_00_19,  
  in_00_21, ou_00_20, in_00_22, ou_00_21, in_00_23, ou_00_22, in_00_24, ou_00_23,  
  in_00_25, ou_00_24;

output 
  in_25_01, ou_25_01, in_25_02, ou_25_02, in_25_03, ou_25_03, in_25_04, ou_25_04,  
  in_25_05, ou_25_05, in_25_06, ou_25_06, in_25_07, ou_25_07, in_25_08, ou_25_08,  
  in_25_09, ou_25_09, in_25_10, ou_25_10, in_25_11, ou_25_11, in_25_12, ou_25_12,  
  in_25_13, ou_25_13, in_25_14, ou_25_14, in_25_15, ou_25_15, in_25_16, ou_25_16,  
  in_25_17, ou_25_17, in_25_18, ou_25_18, in_25_19, ou_25_19, in_25_20, ou_25_20,  
  in_25_21, ou_25_21, in_25_22, ou_25_22, in_25_23, ou_25_23, in_25_24, ou_25_24,  
  in_25_25, ou_25_25;
  wire in_00_01; 
  wire in_00_02; 
  wire in_00_03; 
  wire in_00_04; 
  wire in_00_05; 
  wire in_00_06; 
  wire in_00_07; 
  wire in_00_08; 
  wire in_00_09; 
  wire in_00_10; 
  wire in_00_11; 
  wire in_00_12; 
  wire in_00_13; 
  wire in_00_14; 
  wire in_00_15; 
  wire in_00_16; 
  wire in_00_17; 
  wire in_00_18; 
  wire in_00_19; 
  wire in_00_20; 
  wire in_00_21; 
  wire in_00_22; 
  wire in_00_23; 
  wire in_00_24; 
  wire in_00_25; 
  wire in_01_01; 
  wire in_01_02; 
  wire in_01_03; 
  wire in_01_04; 
  wire in_01_05; 
  wire in_01_06; 
  wire in_01_07; 
  wire in_01_08; 
  wire in_01_09; 
  wire in_01_10; 
  wire in_01_11; 
  wire in_01_12; 
  wire in_01_13; 
  wire in_01_14; 
  wire in_01_15; 
  wire in_01_16; 
  wire in_01_17; 
  wire in_01_18; 
  wire in_01_19; 
  wire in_01_20; 
  wire in_01_21; 
  wire in_01_22; 
  wire in_01_23; 
  wire in_01_24; 
  wire in_01_25; 
  wire in_02_01; 
  wire in_02_02; 
  wire in_02_03; 
  wire in_02_04; 
  wire in_02_05; 
  wire in_02_06; 
  wire in_02_07; 
  wire in_02_08; 
  wire in_02_09; 
  wire in_02_10; 
  wire in_02_11; 
  wire in_02_12; 
  wire in_02_13; 
  wire in_02_14; 
  wire in_02_15; 
  wire in_02_16; 
  wire in_02_17; 
  wire in_02_18; 
  wire in_02_19; 
  wire in_02_20; 
  wire in_02_21; 
  wire in_02_22; 
  wire in_02_23; 
  wire in_02_24; 
  wire in_02_25; 
  wire in_03_01; 
  wire in_03_02; 
  wire in_03_03; 
  wire in_03_04; 
  wire in_03_05; 
  wire in_03_06; 
  wire in_03_07; 
  wire in_03_08; 
  wire in_03_09; 
  wire in_03_10; 
  wire in_03_11; 
  wire in_03_12; 
  wire in_03_13; 
  wire in_03_14; 
  wire in_03_15; 
  wire in_03_16; 
  wire in_03_17; 
  wire in_03_18; 
  wire in_03_19; 
  wire in_03_20; 
  wire in_03_21; 
  wire in_03_22; 
  wire in_03_23; 
  wire in_03_24; 
  wire in_03_25; 
  wire in_04_01; 
  wire in_04_02; 
  wire in_04_03; 
  wire in_04_04; 
  wire in_04_05; 
  wire in_04_06; 
  wire in_04_07; 
  wire in_04_08; 
  wire in_04_09; 
  wire in_04_10; 
  wire in_04_11; 
  wire in_04_12; 
  wire in_04_13; 
  wire in_04_14; 
  wire in_04_15; 
  wire in_04_16; 
  wire in_04_17; 
  wire in_04_18; 
  wire in_04_19; 
  wire in_04_20; 
  wire in_04_21; 
  wire in_04_22; 
  wire in_04_23; 
  wire in_04_24; 
  wire in_04_25; 
  wire in_05_01; 
  wire in_05_02; 
  wire in_05_03; 
  wire in_05_04; 
  wire in_05_05; 
  wire in_05_06; 
  wire in_05_07; 
  wire in_05_08; 
  wire in_05_09; 
  wire in_05_10; 
  wire in_05_11; 
  wire in_05_12; 
  wire in_05_13; 
  wire in_05_14; 
  wire in_05_15; 
  wire in_05_16; 
  wire in_05_17; 
  wire in_05_18; 
  wire in_05_19; 
  wire in_05_20; 
  wire in_05_21; 
  wire in_05_22; 
  wire in_05_23; 
  wire in_05_24; 
  wire in_05_25; 
  wire in_06_01; 
  wire in_06_02; 
  wire in_06_03; 
  wire in_06_04; 
  wire in_06_05; 
  wire in_06_06; 
  wire in_06_07; 
  wire in_06_08; 
  wire in_06_09; 
  wire in_06_10; 
  wire in_06_11; 
  wire in_06_12; 
  wire in_06_13; 
  wire in_06_14; 
  wire in_06_15; 
  wire in_06_16; 
  wire in_06_17; 
  wire in_06_18; 
  wire in_06_19; 
  wire in_06_20; 
  wire in_06_21; 
  wire in_06_22; 
  wire in_06_23; 
  wire in_06_24; 
  wire in_06_25; 
  wire in_07_01; 
  wire in_07_02; 
  wire in_07_03; 
  wire in_07_04; 
  wire in_07_05; 
  wire in_07_06; 
  wire in_07_07; 
  wire in_07_08; 
  wire in_07_09; 
  wire in_07_10; 
  wire in_07_11; 
  wire in_07_12; 
  wire in_07_13; 
  wire in_07_14; 
  wire in_07_15; 
  wire in_07_16; 
  wire in_07_17; 
  wire in_07_18; 
  wire in_07_19; 
  wire in_07_20; 
  wire in_07_21; 
  wire in_07_22; 
  wire in_07_23; 
  wire in_07_24; 
  wire in_07_25; 
  wire in_08_01; 
  wire in_08_02; 
  wire in_08_03; 
  wire in_08_04; 
  wire in_08_05; 
  wire in_08_06; 
  wire in_08_07; 
  wire in_08_08; 
  wire in_08_09; 
  wire in_08_10; 
  wire in_08_11; 
  wire in_08_12; 
  wire in_08_13; 
  wire in_08_14; 
  wire in_08_15; 
  wire in_08_16; 
  wire in_08_17; 
  wire in_08_18; 
  wire in_08_19; 
  wire in_08_20; 
  wire in_08_21; 
  wire in_08_22; 
  wire in_08_23; 
  wire in_08_24; 
  wire in_08_25; 
  wire in_09_01; 
  wire in_09_02; 
  wire in_09_03; 
  wire in_09_04; 
  wire in_09_05; 
  wire in_09_06; 
  wire in_09_07; 
  wire in_09_08; 
  wire in_09_09; 
  wire in_09_10; 
  wire in_09_11; 
  wire in_09_12; 
  wire in_09_13; 
  wire in_09_14; 
  wire in_09_15; 
  wire in_09_16; 
  wire in_09_17; 
  wire in_09_18; 
  wire in_09_19; 
  wire in_09_20; 
  wire in_09_21; 
  wire in_09_22; 
  wire in_09_23; 
  wire in_09_24; 
  wire in_09_25; 
  wire in_10_01; 
  wire in_10_02; 
  wire in_10_03; 
  wire in_10_04; 
  wire in_10_05; 
  wire in_10_06; 
  wire in_10_07; 
  wire in_10_08; 
  wire in_10_09; 
  wire in_10_10; 
  wire in_10_11; 
  wire in_10_12; 
  wire in_10_13; 
  wire in_10_14; 
  wire in_10_15; 
  wire in_10_16; 
  wire in_10_17; 
  wire in_10_18; 
  wire in_10_19; 
  wire in_10_20; 
  wire in_10_21; 
  wire in_10_22; 
  wire in_10_23; 
  wire in_10_24; 
  wire in_10_25; 
  wire in_11_01; 
  wire in_11_02; 
  wire in_11_03; 
  wire in_11_04; 
  wire in_11_05; 
  wire in_11_06; 
  wire in_11_07; 
  wire in_11_08; 
  wire in_11_09; 
  wire in_11_10; 
  wire in_11_11; 
  wire in_11_12; 
  wire in_11_13; 
  wire in_11_14; 
  wire in_11_15; 
  wire in_11_16; 
  wire in_11_17; 
  wire in_11_18; 
  wire in_11_19; 
  wire in_11_20; 
  wire in_11_21; 
  wire in_11_22; 
  wire in_11_23; 
  wire in_11_24; 
  wire in_11_25; 
  wire in_12_01; 
  wire in_12_02; 
  wire in_12_03; 
  wire in_12_04; 
  wire in_12_05; 
  wire in_12_06; 
  wire in_12_07; 
  wire in_12_08; 
  wire in_12_09; 
  wire in_12_10; 
  wire in_12_11; 
  wire in_12_12; 
  wire in_12_13; 
  wire in_12_14; 
  wire in_12_15; 
  wire in_12_16; 
  wire in_12_17; 
  wire in_12_18; 
  wire in_12_19; 
  wire in_12_20; 
  wire in_12_21; 
  wire in_12_22; 
  wire in_12_23; 
  wire in_12_24; 
  wire in_12_25; 
  wire in_13_01; 
  wire in_13_02; 
  wire in_13_03; 
  wire in_13_04; 
  wire in_13_05; 
  wire in_13_06; 
  wire in_13_07; 
  wire in_13_08; 
  wire in_13_09; 
  wire in_13_10; 
  wire in_13_11; 
  wire in_13_12; 
  wire in_13_13; 
  wire in_13_14; 
  wire in_13_15; 
  wire in_13_16; 
  wire in_13_17; 
  wire in_13_18; 
  wire in_13_19; 
  wire in_13_20; 
  wire in_13_21; 
  wire in_13_22; 
  wire in_13_23; 
  wire in_13_24; 
  wire in_13_25; 
  wire in_14_01; 
  wire in_14_02; 
  wire in_14_03; 
  wire in_14_04; 
  wire in_14_05; 
  wire in_14_06; 
  wire in_14_07; 
  wire in_14_08; 
  wire in_14_09; 
  wire in_14_10; 
  wire in_14_11; 
  wire in_14_12; 
  wire in_14_13; 
  wire in_14_14; 
  wire in_14_15; 
  wire in_14_16; 
  wire in_14_17; 
  wire in_14_18; 
  wire in_14_19; 
  wire in_14_20; 
  wire in_14_21; 
  wire in_14_22; 
  wire in_14_23; 
  wire in_14_24; 
  wire in_14_25; 
  wire in_15_01; 
  wire in_15_02; 
  wire in_15_03; 
  wire in_15_04; 
  wire in_15_05; 
  wire in_15_06; 
  wire in_15_07; 
  wire in_15_08; 
  wire in_15_09; 
  wire in_15_10; 
  wire in_15_11; 
  wire in_15_12; 
  wire in_15_13; 
  wire in_15_14; 
  wire in_15_15; 
  wire in_15_16; 
  wire in_15_17; 
  wire in_15_18; 
  wire in_15_19; 
  wire in_15_20; 
  wire in_15_21; 
  wire in_15_22; 
  wire in_15_23; 
  wire in_15_24; 
  wire in_15_25; 
  wire in_16_01; 
  wire in_16_02; 
  wire in_16_03; 
  wire in_16_04; 
  wire in_16_05; 
  wire in_16_06; 
  wire in_16_07; 
  wire in_16_08; 
  wire in_16_09; 
  wire in_16_10; 
  wire in_16_11; 
  wire in_16_12; 
  wire in_16_13; 
  wire in_16_14; 
  wire in_16_15; 
  wire in_16_16; 
  wire in_16_17; 
  wire in_16_18; 
  wire in_16_19; 
  wire in_16_20; 
  wire in_16_21; 
  wire in_16_22; 
  wire in_16_23; 
  wire in_16_24; 
  wire in_16_25; 
  wire in_17_01; 
  wire in_17_02; 
  wire in_17_03; 
  wire in_17_04; 
  wire in_17_05; 
  wire in_17_06; 
  wire in_17_07; 
  wire in_17_08; 
  wire in_17_09; 
  wire in_17_10; 
  wire in_17_11; 
  wire in_17_12; 
  wire in_17_13; 
  wire in_17_14; 
  wire in_17_15; 
  wire in_17_16; 
  wire in_17_17; 
  wire in_17_18; 
  wire in_17_19; 
  wire in_17_20; 
  wire in_17_21; 
  wire in_17_22; 
  wire in_17_23; 
  wire in_17_24; 
  wire in_17_25; 
  wire in_18_01; 
  wire in_18_02; 
  wire in_18_03; 
  wire in_18_04; 
  wire in_18_05; 
  wire in_18_06; 
  wire in_18_07; 
  wire in_18_08; 
  wire in_18_09; 
  wire in_18_10; 
  wire in_18_11; 
  wire in_18_12; 
  wire in_18_13; 
  wire in_18_14; 
  wire in_18_15; 
  wire in_18_16; 
  wire in_18_17; 
  wire in_18_18; 
  wire in_18_19; 
  wire in_18_20; 
  wire in_18_21; 
  wire in_18_22; 
  wire in_18_23; 
  wire in_18_24; 
  wire in_18_25; 
  wire in_19_01; 
  wire in_19_02; 
  wire in_19_03; 
  wire in_19_04; 
  wire in_19_05; 
  wire in_19_06; 
  wire in_19_07; 
  wire in_19_08; 
  wire in_19_09; 
  wire in_19_10; 
  wire in_19_11; 
  wire in_19_12; 
  wire in_19_13; 
  wire in_19_14; 
  wire in_19_15; 
  wire in_19_16; 
  wire in_19_17; 
  wire in_19_18; 
  wire in_19_19; 
  wire in_19_20; 
  wire in_19_21; 
  wire in_19_22; 
  wire in_19_23; 
  wire in_19_24; 
  wire in_19_25; 
  wire in_20_01; 
  wire in_20_02; 
  wire in_20_03; 
  wire in_20_04; 
  wire in_20_05; 
  wire in_20_06; 
  wire in_20_07; 
  wire in_20_08; 
  wire in_20_09; 
  wire in_20_10; 
  wire in_20_11; 
  wire in_20_12; 
  wire in_20_13; 
  wire in_20_14; 
  wire in_20_15; 
  wire in_20_16; 
  wire in_20_17; 
  wire in_20_18; 
  wire in_20_19; 
  wire in_20_20; 
  wire in_20_21; 
  wire in_20_22; 
  wire in_20_23; 
  wire in_20_24; 
  wire in_20_25; 
  wire in_21_01; 
  wire in_21_02; 
  wire in_21_03; 
  wire in_21_04; 
  wire in_21_05; 
  wire in_21_06; 
  wire in_21_07; 
  wire in_21_08; 
  wire in_21_09; 
  wire in_21_10; 
  wire in_21_11; 
  wire in_21_12; 
  wire in_21_13; 
  wire in_21_14; 
  wire in_21_15; 
  wire in_21_16; 
  wire in_21_17; 
  wire in_21_18; 
  wire in_21_19; 
  wire in_21_20; 
  wire in_21_21; 
  wire in_21_22; 
  wire in_21_23; 
  wire in_21_24; 
  wire in_21_25; 
  wire in_22_01; 
  wire in_22_02; 
  wire in_22_03; 
  wire in_22_04; 
  wire in_22_05; 
  wire in_22_06; 
  wire in_22_07; 
  wire in_22_08; 
  wire in_22_09; 
  wire in_22_10; 
  wire in_22_11; 
  wire in_22_12; 
  wire in_22_13; 
  wire in_22_14; 
  wire in_22_15; 
  wire in_22_16; 
  wire in_22_17; 
  wire in_22_18; 
  wire in_22_19; 
  wire in_22_20; 
  wire in_22_21; 
  wire in_22_22; 
  wire in_22_23; 
  wire in_22_24; 
  wire in_22_25; 
  wire in_23_01; 
  wire in_23_02; 
  wire in_23_03; 
  wire in_23_04; 
  wire in_23_05; 
  wire in_23_06; 
  wire in_23_07; 
  wire in_23_08; 
  wire in_23_09; 
  wire in_23_10; 
  wire in_23_11; 
  wire in_23_12; 
  wire in_23_13; 
  wire in_23_14; 
  wire in_23_15; 
  wire in_23_16; 
  wire in_23_17; 
  wire in_23_18; 
  wire in_23_19; 
  wire in_23_20; 
  wire in_23_21; 
  wire in_23_22; 
  wire in_23_23; 
  wire in_23_24; 
  wire in_23_25; 
  wire in_24_01; 
  wire in_24_02; 
  wire in_24_03; 
  wire in_24_04; 
  wire in_24_05; 
  wire in_24_06; 
  wire in_24_07; 
  wire in_24_08; 
  wire in_24_09; 
  wire in_24_10; 
  wire in_24_11; 
  wire in_24_12; 
  wire in_24_13; 
  wire in_24_14; 
  wire in_24_15; 
  wire in_24_16; 
  wire in_24_17; 
  wire in_24_18; 
  wire in_24_19; 
  wire in_24_20; 
  wire in_24_21; 
  wire in_24_22; 
  wire in_24_23; 
  wire in_24_24; 
  wire in_24_25; 

// Instances
  u   u_01_01( clock,enable,reset,set,in_00_01, ou_00_00, in_01_01, ou_01_01 );
  u   u_01_02( clock,enable,reset,set,in_00_02, ou_00_01, in_01_02, ou_01_02 );
  u   u_01_03( clock,enable,reset,set,in_00_03, ou_00_02, in_01_03, ou_01_03 );
  u   u_01_04( clock,enable,reset,set,in_00_04, ou_00_03, in_01_04, ou_01_04 );
  u   u_01_05( clock,enable,reset,set,in_00_05, ou_00_04, in_01_05, ou_01_05 );
  u   u_01_06( clock,enable,reset,set,in_00_06, ou_00_05, in_01_06, ou_01_06 );
  u   u_01_07( clock,enable,reset,set,in_00_07, ou_00_06, in_01_07, ou_01_07 );
  u   u_01_08( clock,enable,reset,set,in_00_08, ou_00_07, in_01_08, ou_01_08 );
  u   u_01_09( clock,enable,reset,set,in_00_09, ou_00_08, in_01_09, ou_01_09 );
  u   u_01_10( clock,enable,reset,set,in_00_10, ou_00_09, in_01_10, ou_01_10 );
  u   u_01_11( clock,enable,reset,set,in_00_11, ou_00_10, in_01_11, ou_01_11 );
  u   u_01_12( clock,enable,reset,set,in_00_12, ou_00_11, in_01_12, ou_01_12 );
  u   u_01_13( clock,enable,reset,set,in_00_13, ou_00_12, in_01_13, ou_01_13 );
  u   u_01_14( clock,enable,reset,set,in_00_14, ou_00_13, in_01_14, ou_01_14 );
  u   u_01_15( clock,enable,reset,set,in_00_15, ou_00_14, in_01_15, ou_01_15 );
  u   u_01_16( clock,enable,reset,set,in_00_16, ou_00_15, in_01_16, ou_01_16 );
  u   u_01_17( clock,enable,reset,set,in_00_17, ou_00_16, in_01_17, ou_01_17 );
  u   u_01_18( clock,enable,reset,set,in_00_18, ou_00_17, in_01_18, ou_01_18 );
  u   u_01_19( clock,enable,reset,set,in_00_19, ou_00_18, in_01_19, ou_01_19 );
  u   u_01_20( clock,enable,reset,set,in_00_20, ou_00_19, in_01_20, ou_01_20 );
  u   u_01_21( clock,enable,reset,set,in_00_21, ou_00_20, in_01_21, ou_01_21 );
  u   u_01_22( clock,enable,reset,set,in_00_22, ou_00_21, in_01_22, ou_01_22 );
  u   u_01_23( clock,enable,reset,set,in_00_23, ou_00_22, in_01_23, ou_01_23 );
  u   u_01_24( clock,enable,reset,set,in_00_24, ou_00_23, in_01_24, ou_01_24 );
  u   u_01_25( clock,enable,reset,set,in_00_25, ou_00_24, in_01_25, ou_01_25 );
  u   u_02_01( clock,enable,reset,set,in_01_01, ou_01_00, in_02_01, ou_02_01 );
  u   u_02_02( clock,enable,reset,set,in_01_02, ou_01_01, in_02_02, ou_02_02 );
  u   u_02_03( clock,enable,reset,set,in_01_03, ou_01_02, in_02_03, ou_02_03 );
  u   u_02_04( clock,enable,reset,set,in_01_04, ou_01_03, in_02_04, ou_02_04 );
  u   u_02_05( clock,enable,reset,set,in_01_05, ou_01_04, in_02_05, ou_02_05 );
  u   u_02_06( clock,enable,reset,set,in_01_06, ou_01_05, in_02_06, ou_02_06 );
  u   u_02_07( clock,enable,reset,set,in_01_07, ou_01_06, in_02_07, ou_02_07 );
  u   u_02_08( clock,enable,reset,set,in_01_08, ou_01_07, in_02_08, ou_02_08 );
  u   u_02_09( clock,enable,reset,set,in_01_09, ou_01_08, in_02_09, ou_02_09 );
  u   u_02_10( clock,enable,reset,set,in_01_10, ou_01_09, in_02_10, ou_02_10 );
  u   u_02_11( clock,enable,reset,set,in_01_11, ou_01_10, in_02_11, ou_02_11 );
  u   u_02_12( clock,enable,reset,set,in_01_12, ou_01_11, in_02_12, ou_02_12 );
  u   u_02_13( clock,enable,reset,set,in_01_13, ou_01_12, in_02_13, ou_02_13 );
  u   u_02_14( clock,enable,reset,set,in_01_14, ou_01_13, in_02_14, ou_02_14 );
  u   u_02_15( clock,enable,reset,set,in_01_15, ou_01_14, in_02_15, ou_02_15 );
  u   u_02_16( clock,enable,reset,set,in_01_16, ou_01_15, in_02_16, ou_02_16 );
  u   u_02_17( clock,enable,reset,set,in_01_17, ou_01_16, in_02_17, ou_02_17 );
  u   u_02_18( clock,enable,reset,set,in_01_18, ou_01_17, in_02_18, ou_02_18 );
  u   u_02_19( clock,enable,reset,set,in_01_19, ou_01_18, in_02_19, ou_02_19 );
  u   u_02_20( clock,enable,reset,set,in_01_20, ou_01_19, in_02_20, ou_02_20 );
  u   u_02_21( clock,enable,reset,set,in_01_21, ou_01_20, in_02_21, ou_02_21 );
  u   u_02_22( clock,enable,reset,set,in_01_22, ou_01_21, in_02_22, ou_02_22 );
  u   u_02_23( clock,enable,reset,set,in_01_23, ou_01_22, in_02_23, ou_02_23 );
  u   u_02_24( clock,enable,reset,set,in_01_24, ou_01_23, in_02_24, ou_02_24 );
  u   u_02_25( clock,enable,reset,set,in_01_25, ou_01_24, in_02_25, ou_02_25 );
  u   u_03_01( clock,enable,reset,set,in_02_01, ou_02_00, in_03_01, ou_03_01 );
  u   u_03_02( clock,enable,reset,set,in_02_02, ou_02_01, in_03_02, ou_03_02 );
  u   u_03_03( clock,enable,reset,set,in_02_03, ou_02_02, in_03_03, ou_03_03 );
  u   u_03_04( clock,enable,reset,set,in_02_04, ou_02_03, in_03_04, ou_03_04 );
  u   u_03_05( clock,enable,reset,set,in_02_05, ou_02_04, in_03_05, ou_03_05 );
  u   u_03_06( clock,enable,reset,set,in_02_06, ou_02_05, in_03_06, ou_03_06 );
  u   u_03_07( clock,enable,reset,set,in_02_07, ou_02_06, in_03_07, ou_03_07 );
  u   u_03_08( clock,enable,reset,set,in_02_08, ou_02_07, in_03_08, ou_03_08 );
  u   u_03_09( clock,enable,reset,set,in_02_09, ou_02_08, in_03_09, ou_03_09 );
  u   u_03_10( clock,enable,reset,set,in_02_10, ou_02_09, in_03_10, ou_03_10 );
  u   u_03_11( clock,enable,reset,set,in_02_11, ou_02_10, in_03_11, ou_03_11 );
  u   u_03_12( clock,enable,reset,set,in_02_12, ou_02_11, in_03_12, ou_03_12 );
  u   u_03_13( clock,enable,reset,set,in_02_13, ou_02_12, in_03_13, ou_03_13 );
  u   u_03_14( clock,enable,reset,set,in_02_14, ou_02_13, in_03_14, ou_03_14 );
  u   u_03_15( clock,enable,reset,set,in_02_15, ou_02_14, in_03_15, ou_03_15 );
  u   u_03_16( clock,enable,reset,set,in_02_16, ou_02_15, in_03_16, ou_03_16 );
  u   u_03_17( clock,enable,reset,set,in_02_17, ou_02_16, in_03_17, ou_03_17 );
  u   u_03_18( clock,enable,reset,set,in_02_18, ou_02_17, in_03_18, ou_03_18 );
  u   u_03_19( clock,enable,reset,set,in_02_19, ou_02_18, in_03_19, ou_03_19 );
  u   u_03_20( clock,enable,reset,set,in_02_20, ou_02_19, in_03_20, ou_03_20 );
  u   u_03_21( clock,enable,reset,set,in_02_21, ou_02_20, in_03_21, ou_03_21 );
  u   u_03_22( clock,enable,reset,set,in_02_22, ou_02_21, in_03_22, ou_03_22 );
  u   u_03_23( clock,enable,reset,set,in_02_23, ou_02_22, in_03_23, ou_03_23 );
  u   u_03_24( clock,enable,reset,set,in_02_24, ou_02_23, in_03_24, ou_03_24 );
  u   u_03_25( clock,enable,reset,set,in_02_25, ou_02_24, in_03_25, ou_03_25 );
  u   u_04_01( clock,enable,reset,set,in_03_01, ou_03_00, in_04_01, ou_04_01 );
  u   u_04_02( clock,enable,reset,set,in_03_02, ou_03_01, in_04_02, ou_04_02 );
  u   u_04_03( clock,enable,reset,set,in_03_03, ou_03_02, in_04_03, ou_04_03 );
  u   u_04_04( clock,enable,reset,set,in_03_04, ou_03_03, in_04_04, ou_04_04 );
  u   u_04_05( clock,enable,reset,set,in_03_05, ou_03_04, in_04_05, ou_04_05 );
  u   u_04_06( clock,enable,reset,set,in_03_06, ou_03_05, in_04_06, ou_04_06 );
  u   u_04_07( clock,enable,reset,set,in_03_07, ou_03_06, in_04_07, ou_04_07 );
  u   u_04_08( clock,enable,reset,set,in_03_08, ou_03_07, in_04_08, ou_04_08 );
  u   u_04_09( clock,enable,reset,set,in_03_09, ou_03_08, in_04_09, ou_04_09 );
  u   u_04_10( clock,enable,reset,set,in_03_10, ou_03_09, in_04_10, ou_04_10 );
  u   u_04_11( clock,enable,reset,set,in_03_11, ou_03_10, in_04_11, ou_04_11 );
  u   u_04_12( clock,enable,reset,set,in_03_12, ou_03_11, in_04_12, ou_04_12 );
  u   u_04_13( clock,enable,reset,set,in_03_13, ou_03_12, in_04_13, ou_04_13 );
  u   u_04_14( clock,enable,reset,set,in_03_14, ou_03_13, in_04_14, ou_04_14 );
  u   u_04_15( clock,enable,reset,set,in_03_15, ou_03_14, in_04_15, ou_04_15 );
  u   u_04_16( clock,enable,reset,set,in_03_16, ou_03_15, in_04_16, ou_04_16 );
  u   u_04_17( clock,enable,reset,set,in_03_17, ou_03_16, in_04_17, ou_04_17 );
  u   u_04_18( clock,enable,reset,set,in_03_18, ou_03_17, in_04_18, ou_04_18 );
  u   u_04_19( clock,enable,reset,set,in_03_19, ou_03_18, in_04_19, ou_04_19 );
  u   u_04_20( clock,enable,reset,set,in_03_20, ou_03_19, in_04_20, ou_04_20 );
  u   u_04_21( clock,enable,reset,set,in_03_21, ou_03_20, in_04_21, ou_04_21 );
  u   u_04_22( clock,enable,reset,set,in_03_22, ou_03_21, in_04_22, ou_04_22 );
  u   u_04_23( clock,enable,reset,set,in_03_23, ou_03_22, in_04_23, ou_04_23 );
  u   u_04_24( clock,enable,reset,set,in_03_24, ou_03_23, in_04_24, ou_04_24 );
  u   u_04_25( clock,enable,reset,set,in_03_25, ou_03_24, in_04_25, ou_04_25 );
  u   u_05_01( clock,enable,reset,set,in_04_01, ou_04_00, in_05_01, ou_05_01 );
  u   u_05_02( clock,enable,reset,set,in_04_02, ou_04_01, in_05_02, ou_05_02 );
  u   u_05_03( clock,enable,reset,set,in_04_03, ou_04_02, in_05_03, ou_05_03 );
  u   u_05_04( clock,enable,reset,set,in_04_04, ou_04_03, in_05_04, ou_05_04 );
  u   u_05_05( clock,enable,reset,set,in_04_05, ou_04_04, in_05_05, ou_05_05 );
  u   u_05_06( clock,enable,reset,set,in_04_06, ou_04_05, in_05_06, ou_05_06 );
  u   u_05_07( clock,enable,reset,set,in_04_07, ou_04_06, in_05_07, ou_05_07 );
  u   u_05_08( clock,enable,reset,set,in_04_08, ou_04_07, in_05_08, ou_05_08 );
  u   u_05_09( clock,enable,reset,set,in_04_09, ou_04_08, in_05_09, ou_05_09 );
  u   u_05_10( clock,enable,reset,set,in_04_10, ou_04_09, in_05_10, ou_05_10 );
  u   u_05_11( clock,enable,reset,set,in_04_11, ou_04_10, in_05_11, ou_05_11 );
  u   u_05_12( clock,enable,reset,set,in_04_12, ou_04_11, in_05_12, ou_05_12 );
  u   u_05_13( clock,enable,reset,set,in_04_13, ou_04_12, in_05_13, ou_05_13 );
  u   u_05_14( clock,enable,reset,set,in_04_14, ou_04_13, in_05_14, ou_05_14 );
  u   u_05_15( clock,enable,reset,set,in_04_15, ou_04_14, in_05_15, ou_05_15 );
  u   u_05_16( clock,enable,reset,set,in_04_16, ou_04_15, in_05_16, ou_05_16 );
  u   u_05_17( clock,enable,reset,set,in_04_17, ou_04_16, in_05_17, ou_05_17 );
  u   u_05_18( clock,enable,reset,set,in_04_18, ou_04_17, in_05_18, ou_05_18 );
  u   u_05_19( clock,enable,reset,set,in_04_19, ou_04_18, in_05_19, ou_05_19 );
  u   u_05_20( clock,enable,reset,set,in_04_20, ou_04_19, in_05_20, ou_05_20 );
  u   u_05_21( clock,enable,reset,set,in_04_21, ou_04_20, in_05_21, ou_05_21 );
  u   u_05_22( clock,enable,reset,set,in_04_22, ou_04_21, in_05_22, ou_05_22 );
  u   u_05_23( clock,enable,reset,set,in_04_23, ou_04_22, in_05_23, ou_05_23 );
  u   u_05_24( clock,enable,reset,set,in_04_24, ou_04_23, in_05_24, ou_05_24 );
  u   u_05_25( clock,enable,reset,set,in_04_25, ou_04_24, in_05_25, ou_05_25 );
  u   u_06_01( clock,enable,reset,set,in_05_01, ou_05_00, in_06_01, ou_06_01 );
  u   u_06_02( clock,enable,reset,set,in_05_02, ou_05_01, in_06_02, ou_06_02 );
  u   u_06_03( clock,enable,reset,set,in_05_03, ou_05_02, in_06_03, ou_06_03 );
  u   u_06_04( clock,enable,reset,set,in_05_04, ou_05_03, in_06_04, ou_06_04 );
  u   u_06_05( clock,enable,reset,set,in_05_05, ou_05_04, in_06_05, ou_06_05 );
  u   u_06_06( clock,enable,reset,set,in_05_06, ou_05_05, in_06_06, ou_06_06 );
  u   u_06_07( clock,enable,reset,set,in_05_07, ou_05_06, in_06_07, ou_06_07 );
  u   u_06_08( clock,enable,reset,set,in_05_08, ou_05_07, in_06_08, ou_06_08 );
  u   u_06_09( clock,enable,reset,set,in_05_09, ou_05_08, in_06_09, ou_06_09 );
  u   u_06_10( clock,enable,reset,set,in_05_10, ou_05_09, in_06_10, ou_06_10 );
  u   u_06_11( clock,enable,reset,set,in_05_11, ou_05_10, in_06_11, ou_06_11 );
  u   u_06_12( clock,enable,reset,set,in_05_12, ou_05_11, in_06_12, ou_06_12 );
  u   u_06_13( clock,enable,reset,set,in_05_13, ou_05_12, in_06_13, ou_06_13 );
  u   u_06_14( clock,enable,reset,set,in_05_14, ou_05_13, in_06_14, ou_06_14 );
  u   u_06_15( clock,enable,reset,set,in_05_15, ou_05_14, in_06_15, ou_06_15 );
  u   u_06_16( clock,enable,reset,set,in_05_16, ou_05_15, in_06_16, ou_06_16 );
  u   u_06_17( clock,enable,reset,set,in_05_17, ou_05_16, in_06_17, ou_06_17 );
  u   u_06_18( clock,enable,reset,set,in_05_18, ou_05_17, in_06_18, ou_06_18 );
  u   u_06_19( clock,enable,reset,set,in_05_19, ou_05_18, in_06_19, ou_06_19 );
  u   u_06_20( clock,enable,reset,set,in_05_20, ou_05_19, in_06_20, ou_06_20 );
  u   u_06_21( clock,enable,reset,set,in_05_21, ou_05_20, in_06_21, ou_06_21 );
  u   u_06_22( clock,enable,reset,set,in_05_22, ou_05_21, in_06_22, ou_06_22 );
  u   u_06_23( clock,enable,reset,set,in_05_23, ou_05_22, in_06_23, ou_06_23 );
  u   u_06_24( clock,enable,reset,set,in_05_24, ou_05_23, in_06_24, ou_06_24 );
  u   u_06_25( clock,enable,reset,set,in_05_25, ou_05_24, in_06_25, ou_06_25 );
  u   u_07_01( clock,enable,reset,set,in_06_01, ou_06_00, in_07_01, ou_07_01 );
  u   u_07_02( clock,enable,reset,set,in_06_02, ou_06_01, in_07_02, ou_07_02 );
  u   u_07_03( clock,enable,reset,set,in_06_03, ou_06_02, in_07_03, ou_07_03 );
  u   u_07_04( clock,enable,reset,set,in_06_04, ou_06_03, in_07_04, ou_07_04 );
  u   u_07_05( clock,enable,reset,set,in_06_05, ou_06_04, in_07_05, ou_07_05 );
  u   u_07_06( clock,enable,reset,set,in_06_06, ou_06_05, in_07_06, ou_07_06 );
  u   u_07_07( clock,enable,reset,set,in_06_07, ou_06_06, in_07_07, ou_07_07 );
  u   u_07_08( clock,enable,reset,set,in_06_08, ou_06_07, in_07_08, ou_07_08 );
  u   u_07_09( clock,enable,reset,set,in_06_09, ou_06_08, in_07_09, ou_07_09 );
  u   u_07_10( clock,enable,reset,set,in_06_10, ou_06_09, in_07_10, ou_07_10 );
  u   u_07_11( clock,enable,reset,set,in_06_11, ou_06_10, in_07_11, ou_07_11 );
  u   u_07_12( clock,enable,reset,set,in_06_12, ou_06_11, in_07_12, ou_07_12 );
  u   u_07_13( clock,enable,reset,set,in_06_13, ou_06_12, in_07_13, ou_07_13 );
  u   u_07_14( clock,enable,reset,set,in_06_14, ou_06_13, in_07_14, ou_07_14 );
  u   u_07_15( clock,enable,reset,set,in_06_15, ou_06_14, in_07_15, ou_07_15 );
  u   u_07_16( clock,enable,reset,set,in_06_16, ou_06_15, in_07_16, ou_07_16 );
  u   u_07_17( clock,enable,reset,set,in_06_17, ou_06_16, in_07_17, ou_07_17 );
  u   u_07_18( clock,enable,reset,set,in_06_18, ou_06_17, in_07_18, ou_07_18 );
  u   u_07_19( clock,enable,reset,set,in_06_19, ou_06_18, in_07_19, ou_07_19 );
  u   u_07_20( clock,enable,reset,set,in_06_20, ou_06_19, in_07_20, ou_07_20 );
  u   u_07_21( clock,enable,reset,set,in_06_21, ou_06_20, in_07_21, ou_07_21 );
  u   u_07_22( clock,enable,reset,set,in_06_22, ou_06_21, in_07_22, ou_07_22 );
  u   u_07_23( clock,enable,reset,set,in_06_23, ou_06_22, in_07_23, ou_07_23 );
  u   u_07_24( clock,enable,reset,set,in_06_24, ou_06_23, in_07_24, ou_07_24 );
  u   u_07_25( clock,enable,reset,set,in_06_25, ou_06_24, in_07_25, ou_07_25 );
  u   u_08_01( clock,enable,reset,set,in_07_01, ou_07_00, in_08_01, ou_08_01 );
  u   u_08_02( clock,enable,reset,set,in_07_02, ou_07_01, in_08_02, ou_08_02 );
  u   u_08_03( clock,enable,reset,set,in_07_03, ou_07_02, in_08_03, ou_08_03 );
  u   u_08_04( clock,enable,reset,set,in_07_04, ou_07_03, in_08_04, ou_08_04 );
  u   u_08_05( clock,enable,reset,set,in_07_05, ou_07_04, in_08_05, ou_08_05 );
  u   u_08_06( clock,enable,reset,set,in_07_06, ou_07_05, in_08_06, ou_08_06 );
  u   u_08_07( clock,enable,reset,set,in_07_07, ou_07_06, in_08_07, ou_08_07 );
  u   u_08_08( clock,enable,reset,set,in_07_08, ou_07_07, in_08_08, ou_08_08 );
  u   u_08_09( clock,enable,reset,set,in_07_09, ou_07_08, in_08_09, ou_08_09 );
  u   u_08_10( clock,enable,reset,set,in_07_10, ou_07_09, in_08_10, ou_08_10 );
  u   u_08_11( clock,enable,reset,set,in_07_11, ou_07_10, in_08_11, ou_08_11 );
  u   u_08_12( clock,enable,reset,set,in_07_12, ou_07_11, in_08_12, ou_08_12 );
  u   u_08_13( clock,enable,reset,set,in_07_13, ou_07_12, in_08_13, ou_08_13 );
  u   u_08_14( clock,enable,reset,set,in_07_14, ou_07_13, in_08_14, ou_08_14 );
  u   u_08_15( clock,enable,reset,set,in_07_15, ou_07_14, in_08_15, ou_08_15 );
  u   u_08_16( clock,enable,reset,set,in_07_16, ou_07_15, in_08_16, ou_08_16 );
  u   u_08_17( clock,enable,reset,set,in_07_17, ou_07_16, in_08_17, ou_08_17 );
  u   u_08_18( clock,enable,reset,set,in_07_18, ou_07_17, in_08_18, ou_08_18 );
  u   u_08_19( clock,enable,reset,set,in_07_19, ou_07_18, in_08_19, ou_08_19 );
  u   u_08_20( clock,enable,reset,set,in_07_20, ou_07_19, in_08_20, ou_08_20 );
  u   u_08_21( clock,enable,reset,set,in_07_21, ou_07_20, in_08_21, ou_08_21 );
  u   u_08_22( clock,enable,reset,set,in_07_22, ou_07_21, in_08_22, ou_08_22 );
  u   u_08_23( clock,enable,reset,set,in_07_23, ou_07_22, in_08_23, ou_08_23 );
  u   u_08_24( clock,enable,reset,set,in_07_24, ou_07_23, in_08_24, ou_08_24 );
  u   u_08_25( clock,enable,reset,set,in_07_25, ou_07_24, in_08_25, ou_08_25 );
  u   u_09_01( clock,enable,reset,set,in_08_01, ou_08_00, in_09_01, ou_09_01 );
  u   u_09_02( clock,enable,reset,set,in_08_02, ou_08_01, in_09_02, ou_09_02 );
  u   u_09_03( clock,enable,reset,set,in_08_03, ou_08_02, in_09_03, ou_09_03 );
  u   u_09_04( clock,enable,reset,set,in_08_04, ou_08_03, in_09_04, ou_09_04 );
  u   u_09_05( clock,enable,reset,set,in_08_05, ou_08_04, in_09_05, ou_09_05 );
  u   u_09_06( clock,enable,reset,set,in_08_06, ou_08_05, in_09_06, ou_09_06 );
  u   u_09_07( clock,enable,reset,set,in_08_07, ou_08_06, in_09_07, ou_09_07 );
  u   u_09_08( clock,enable,reset,set,in_08_08, ou_08_07, in_09_08, ou_09_08 );
  u   u_09_09( clock,enable,reset,set,in_08_09, ou_08_08, in_09_09, ou_09_09 );
  u   u_09_10( clock,enable,reset,set,in_08_10, ou_08_09, in_09_10, ou_09_10 );
  u   u_09_11( clock,enable,reset,set,in_08_11, ou_08_10, in_09_11, ou_09_11 );
  u   u_09_12( clock,enable,reset,set,in_08_12, ou_08_11, in_09_12, ou_09_12 );
  u   u_09_13( clock,enable,reset,set,in_08_13, ou_08_12, in_09_13, ou_09_13 );
  u   u_09_14( clock,enable,reset,set,in_08_14, ou_08_13, in_09_14, ou_09_14 );
  u   u_09_15( clock,enable,reset,set,in_08_15, ou_08_14, in_09_15, ou_09_15 );
  u   u_09_16( clock,enable,reset,set,in_08_16, ou_08_15, in_09_16, ou_09_16 );
  u   u_09_17( clock,enable,reset,set,in_08_17, ou_08_16, in_09_17, ou_09_17 );
  u   u_09_18( clock,enable,reset,set,in_08_18, ou_08_17, in_09_18, ou_09_18 );
  u   u_09_19( clock,enable,reset,set,in_08_19, ou_08_18, in_09_19, ou_09_19 );
  u   u_09_20( clock,enable,reset,set,in_08_20, ou_08_19, in_09_20, ou_09_20 );
  u   u_09_21( clock,enable,reset,set,in_08_21, ou_08_20, in_09_21, ou_09_21 );
  u   u_09_22( clock,enable,reset,set,in_08_22, ou_08_21, in_09_22, ou_09_22 );
  u   u_09_23( clock,enable,reset,set,in_08_23, ou_08_22, in_09_23, ou_09_23 );
  u   u_09_24( clock,enable,reset,set,in_08_24, ou_08_23, in_09_24, ou_09_24 );
  u   u_09_25( clock,enable,reset,set,in_08_25, ou_08_24, in_09_25, ou_09_25 );
  u   u_10_01( clock,enable,reset,set,in_09_01, ou_09_00, in_10_01, ou_10_01 );
  u   u_10_02( clock,enable,reset,set,in_09_02, ou_09_01, in_10_02, ou_10_02 );
  u   u_10_03( clock,enable,reset,set,in_09_03, ou_09_02, in_10_03, ou_10_03 );
  u   u_10_04( clock,enable,reset,set,in_09_04, ou_09_03, in_10_04, ou_10_04 );
  u   u_10_05( clock,enable,reset,set,in_09_05, ou_09_04, in_10_05, ou_10_05 );
  u   u_10_06( clock,enable,reset,set,in_09_06, ou_09_05, in_10_06, ou_10_06 );
  u   u_10_07( clock,enable,reset,set,in_09_07, ou_09_06, in_10_07, ou_10_07 );
  u   u_10_08( clock,enable,reset,set,in_09_08, ou_09_07, in_10_08, ou_10_08 );
  u   u_10_09( clock,enable,reset,set,in_09_09, ou_09_08, in_10_09, ou_10_09 );
  u   u_10_10( clock,enable,reset,set,in_09_10, ou_09_09, in_10_10, ou_10_10 );
  u   u_10_11( clock,enable,reset,set,in_09_11, ou_09_10, in_10_11, ou_10_11 );
  u   u_10_12( clock,enable,reset,set,in_09_12, ou_09_11, in_10_12, ou_10_12 );
  u   u_10_13( clock,enable,reset,set,in_09_13, ou_09_12, in_10_13, ou_10_13 );
  u   u_10_14( clock,enable,reset,set,in_09_14, ou_09_13, in_10_14, ou_10_14 );
  u   u_10_15( clock,enable,reset,set,in_09_15, ou_09_14, in_10_15, ou_10_15 );
  u   u_10_16( clock,enable,reset,set,in_09_16, ou_09_15, in_10_16, ou_10_16 );
  u   u_10_17( clock,enable,reset,set,in_09_17, ou_09_16, in_10_17, ou_10_17 );
  u   u_10_18( clock,enable,reset,set,in_09_18, ou_09_17, in_10_18, ou_10_18 );
  u   u_10_19( clock,enable,reset,set,in_09_19, ou_09_18, in_10_19, ou_10_19 );
  u   u_10_20( clock,enable,reset,set,in_09_20, ou_09_19, in_10_20, ou_10_20 );
  u   u_10_21( clock,enable,reset,set,in_09_21, ou_09_20, in_10_21, ou_10_21 );
  u   u_10_22( clock,enable,reset,set,in_09_22, ou_09_21, in_10_22, ou_10_22 );
  u   u_10_23( clock,enable,reset,set,in_09_23, ou_09_22, in_10_23, ou_10_23 );
  u   u_10_24( clock,enable,reset,set,in_09_24, ou_09_23, in_10_24, ou_10_24 );
  u   u_10_25( clock,enable,reset,set,in_09_25, ou_09_24, in_10_25, ou_10_25 );
  u   u_11_01( clock,enable,reset,set,in_10_01, ou_10_00, in_11_01, ou_11_01 );
  u   u_11_02( clock,enable,reset,set,in_10_02, ou_10_01, in_11_02, ou_11_02 );
  u   u_11_03( clock,enable,reset,set,in_10_03, ou_10_02, in_11_03, ou_11_03 );
  u   u_11_04( clock,enable,reset,set,in_10_04, ou_10_03, in_11_04, ou_11_04 );
  u   u_11_05( clock,enable,reset,set,in_10_05, ou_10_04, in_11_05, ou_11_05 );
  u   u_11_06( clock,enable,reset,set,in_10_06, ou_10_05, in_11_06, ou_11_06 );
  u   u_11_07( clock,enable,reset,set,in_10_07, ou_10_06, in_11_07, ou_11_07 );
  u   u_11_08( clock,enable,reset,set,in_10_08, ou_10_07, in_11_08, ou_11_08 );
  u   u_11_09( clock,enable,reset,set,in_10_09, ou_10_08, in_11_09, ou_11_09 );
  u   u_11_10( clock,enable,reset,set,in_10_10, ou_10_09, in_11_10, ou_11_10 );
  u   u_11_11( clock,enable,reset,set,in_10_11, ou_10_10, in_11_11, ou_11_11 );
  u   u_11_12( clock,enable,reset,set,in_10_12, ou_10_11, in_11_12, ou_11_12 );
  u   u_11_13( clock,enable,reset,set,in_10_13, ou_10_12, in_11_13, ou_11_13 );
  u   u_11_14( clock,enable,reset,set,in_10_14, ou_10_13, in_11_14, ou_11_14 );
  u   u_11_15( clock,enable,reset,set,in_10_15, ou_10_14, in_11_15, ou_11_15 );
  u   u_11_16( clock,enable,reset,set,in_10_16, ou_10_15, in_11_16, ou_11_16 );
  u   u_11_17( clock,enable,reset,set,in_10_17, ou_10_16, in_11_17, ou_11_17 );
  u   u_11_18( clock,enable,reset,set,in_10_18, ou_10_17, in_11_18, ou_11_18 );
  u   u_11_19( clock,enable,reset,set,in_10_19, ou_10_18, in_11_19, ou_11_19 );
  u   u_11_20( clock,enable,reset,set,in_10_20, ou_10_19, in_11_20, ou_11_20 );
  u   u_11_21( clock,enable,reset,set,in_10_21, ou_10_20, in_11_21, ou_11_21 );
  u   u_11_22( clock,enable,reset,set,in_10_22, ou_10_21, in_11_22, ou_11_22 );
  u   u_11_23( clock,enable,reset,set,in_10_23, ou_10_22, in_11_23, ou_11_23 );
  u   u_11_24( clock,enable,reset,set,in_10_24, ou_10_23, in_11_24, ou_11_24 );
  u   u_11_25( clock,enable,reset,set,in_10_25, ou_10_24, in_11_25, ou_11_25 );
  u   u_12_01( clock,enable,reset,set,in_11_01, ou_11_00, in_12_01, ou_12_01 );
  u   u_12_02( clock,enable,reset,set,in_11_02, ou_11_01, in_12_02, ou_12_02 );
  u   u_12_03( clock,enable,reset,set,in_11_03, ou_11_02, in_12_03, ou_12_03 );
  u   u_12_04( clock,enable,reset,set,in_11_04, ou_11_03, in_12_04, ou_12_04 );
  u   u_12_05( clock,enable,reset,set,in_11_05, ou_11_04, in_12_05, ou_12_05 );
  u   u_12_06( clock,enable,reset,set,in_11_06, ou_11_05, in_12_06, ou_12_06 );
  u   u_12_07( clock,enable,reset,set,in_11_07, ou_11_06, in_12_07, ou_12_07 );
  u   u_12_08( clock,enable,reset,set,in_11_08, ou_11_07, in_12_08, ou_12_08 );
  u   u_12_09( clock,enable,reset,set,in_11_09, ou_11_08, in_12_09, ou_12_09 );
  u   u_12_10( clock,enable,reset,set,in_11_10, ou_11_09, in_12_10, ou_12_10 );
  u   u_12_11( clock,enable,reset,set,in_11_11, ou_11_10, in_12_11, ou_12_11 );
  u   u_12_12( clock,enable,reset,set,in_11_12, ou_11_11, in_12_12, ou_12_12 );
  u   u_12_13( clock,enable,reset,set,in_11_13, ou_11_12, in_12_13, ou_12_13 );
  u   u_12_14( clock,enable,reset,set,in_11_14, ou_11_13, in_12_14, ou_12_14 );
  u   u_12_15( clock,enable,reset,set,in_11_15, ou_11_14, in_12_15, ou_12_15 );
  u   u_12_16( clock,enable,reset,set,in_11_16, ou_11_15, in_12_16, ou_12_16 );
  u   u_12_17( clock,enable,reset,set,in_11_17, ou_11_16, in_12_17, ou_12_17 );
  u   u_12_18( clock,enable,reset,set,in_11_18, ou_11_17, in_12_18, ou_12_18 );
  u   u_12_19( clock,enable,reset,set,in_11_19, ou_11_18, in_12_19, ou_12_19 );
  u   u_12_20( clock,enable,reset,set,in_11_20, ou_11_19, in_12_20, ou_12_20 );
  u   u_12_21( clock,enable,reset,set,in_11_21, ou_11_20, in_12_21, ou_12_21 );
  u   u_12_22( clock,enable,reset,set,in_11_22, ou_11_21, in_12_22, ou_12_22 );
  u   u_12_23( clock,enable,reset,set,in_11_23, ou_11_22, in_12_23, ou_12_23 );
  u   u_12_24( clock,enable,reset,set,in_11_24, ou_11_23, in_12_24, ou_12_24 );
  u   u_12_25( clock,enable,reset,set,in_11_25, ou_11_24, in_12_25, ou_12_25 );
  u   u_13_01( clock,enable,reset,set,in_12_01, ou_12_00, in_13_01, ou_13_01 );
  u   u_13_02( clock,enable,reset,set,in_12_02, ou_12_01, in_13_02, ou_13_02 );
  u   u_13_03( clock,enable,reset,set,in_12_03, ou_12_02, in_13_03, ou_13_03 );
  u   u_13_04( clock,enable,reset,set,in_12_04, ou_12_03, in_13_04, ou_13_04 );
  u   u_13_05( clock,enable,reset,set,in_12_05, ou_12_04, in_13_05, ou_13_05 );
  u   u_13_06( clock,enable,reset,set,in_12_06, ou_12_05, in_13_06, ou_13_06 );
  u   u_13_07( clock,enable,reset,set,in_12_07, ou_12_06, in_13_07, ou_13_07 );
  u   u_13_08( clock,enable,reset,set,in_12_08, ou_12_07, in_13_08, ou_13_08 );
  u   u_13_09( clock,enable,reset,set,in_12_09, ou_12_08, in_13_09, ou_13_09 );
  u   u_13_10( clock,enable,reset,set,in_12_10, ou_12_09, in_13_10, ou_13_10 );
  u   u_13_11( clock,enable,reset,set,in_12_11, ou_12_10, in_13_11, ou_13_11 );
  u   u_13_12( clock,enable,reset,set,in_12_12, ou_12_11, in_13_12, ou_13_12 );
  u   u_13_13( clock,enable,reset,set,in_12_13, ou_12_12, in_13_13, ou_13_13 );
  u   u_13_14( clock,enable,reset,set,in_12_14, ou_12_13, in_13_14, ou_13_14 );
  u   u_13_15( clock,enable,reset,set,in_12_15, ou_12_14, in_13_15, ou_13_15 );
  u   u_13_16( clock,enable,reset,set,in_12_16, ou_12_15, in_13_16, ou_13_16 );
  u   u_13_17( clock,enable,reset,set,in_12_17, ou_12_16, in_13_17, ou_13_17 );
  u   u_13_18( clock,enable,reset,set,in_12_18, ou_12_17, in_13_18, ou_13_18 );
  u   u_13_19( clock,enable,reset,set,in_12_19, ou_12_18, in_13_19, ou_13_19 );
  u   u_13_20( clock,enable,reset,set,in_12_20, ou_12_19, in_13_20, ou_13_20 );
  u   u_13_21( clock,enable,reset,set,in_12_21, ou_12_20, in_13_21, ou_13_21 );
  u   u_13_22( clock,enable,reset,set,in_12_22, ou_12_21, in_13_22, ou_13_22 );
  u   u_13_23( clock,enable,reset,set,in_12_23, ou_12_22, in_13_23, ou_13_23 );
  u   u_13_24( clock,enable,reset,set,in_12_24, ou_12_23, in_13_24, ou_13_24 );
  u   u_13_25( clock,enable,reset,set,in_12_25, ou_12_24, in_13_25, ou_13_25 );
  u   u_14_01( clock,enable,reset,set,in_13_01, ou_13_00, in_14_01, ou_14_01 );
  u   u_14_02( clock,enable,reset,set,in_13_02, ou_13_01, in_14_02, ou_14_02 );
  u   u_14_03( clock,enable,reset,set,in_13_03, ou_13_02, in_14_03, ou_14_03 );
  u   u_14_04( clock,enable,reset,set,in_13_04, ou_13_03, in_14_04, ou_14_04 );
  u   u_14_05( clock,enable,reset,set,in_13_05, ou_13_04, in_14_05, ou_14_05 );
  u   u_14_06( clock,enable,reset,set,in_13_06, ou_13_05, in_14_06, ou_14_06 );
  u   u_14_07( clock,enable,reset,set,in_13_07, ou_13_06, in_14_07, ou_14_07 );
  u   u_14_08( clock,enable,reset,set,in_13_08, ou_13_07, in_14_08, ou_14_08 );
  u   u_14_09( clock,enable,reset,set,in_13_09, ou_13_08, in_14_09, ou_14_09 );
  u   u_14_10( clock,enable,reset,set,in_13_10, ou_13_09, in_14_10, ou_14_10 );
  u   u_14_11( clock,enable,reset,set,in_13_11, ou_13_10, in_14_11, ou_14_11 );
  u   u_14_12( clock,enable,reset,set,in_13_12, ou_13_11, in_14_12, ou_14_12 );
  u   u_14_13( clock,enable,reset,set,in_13_13, ou_13_12, in_14_13, ou_14_13 );
  u   u_14_14( clock,enable,reset,set,in_13_14, ou_13_13, in_14_14, ou_14_14 );
  u   u_14_15( clock,enable,reset,set,in_13_15, ou_13_14, in_14_15, ou_14_15 );
  u   u_14_16( clock,enable,reset,set,in_13_16, ou_13_15, in_14_16, ou_14_16 );
  u   u_14_17( clock,enable,reset,set,in_13_17, ou_13_16, in_14_17, ou_14_17 );
  u   u_14_18( clock,enable,reset,set,in_13_18, ou_13_17, in_14_18, ou_14_18 );
  u   u_14_19( clock,enable,reset,set,in_13_19, ou_13_18, in_14_19, ou_14_19 );
  u   u_14_20( clock,enable,reset,set,in_13_20, ou_13_19, in_14_20, ou_14_20 );
  u   u_14_21( clock,enable,reset,set,in_13_21, ou_13_20, in_14_21, ou_14_21 );
  u   u_14_22( clock,enable,reset,set,in_13_22, ou_13_21, in_14_22, ou_14_22 );
  u   u_14_23( clock,enable,reset,set,in_13_23, ou_13_22, in_14_23, ou_14_23 );
  u   u_14_24( clock,enable,reset,set,in_13_24, ou_13_23, in_14_24, ou_14_24 );
  u   u_14_25( clock,enable,reset,set,in_13_25, ou_13_24, in_14_25, ou_14_25 );
  u   u_15_01( clock,enable,reset,set,in_14_01, ou_14_00, in_15_01, ou_15_01 );
  u   u_15_02( clock,enable,reset,set,in_14_02, ou_14_01, in_15_02, ou_15_02 );
  u   u_15_03( clock,enable,reset,set,in_14_03, ou_14_02, in_15_03, ou_15_03 );
  u   u_15_04( clock,enable,reset,set,in_14_04, ou_14_03, in_15_04, ou_15_04 );
  u   u_15_05( clock,enable,reset,set,in_14_05, ou_14_04, in_15_05, ou_15_05 );
  u   u_15_06( clock,enable,reset,set,in_14_06, ou_14_05, in_15_06, ou_15_06 );
  u   u_15_07( clock,enable,reset,set,in_14_07, ou_14_06, in_15_07, ou_15_07 );
  u   u_15_08( clock,enable,reset,set,in_14_08, ou_14_07, in_15_08, ou_15_08 );
  u   u_15_09( clock,enable,reset,set,in_14_09, ou_14_08, in_15_09, ou_15_09 );
  u   u_15_10( clock,enable,reset,set,in_14_10, ou_14_09, in_15_10, ou_15_10 );
  u   u_15_11( clock,enable,reset,set,in_14_11, ou_14_10, in_15_11, ou_15_11 );
  u   u_15_12( clock,enable,reset,set,in_14_12, ou_14_11, in_15_12, ou_15_12 );
  u   u_15_13( clock,enable,reset,set,in_14_13, ou_14_12, in_15_13, ou_15_13 );
  u   u_15_14( clock,enable,reset,set,in_14_14, ou_14_13, in_15_14, ou_15_14 );
  u   u_15_15( clock,enable,reset,set,in_14_15, ou_14_14, in_15_15, ou_15_15 );
  u   u_15_16( clock,enable,reset,set,in_14_16, ou_14_15, in_15_16, ou_15_16 );
  u   u_15_17( clock,enable,reset,set,in_14_17, ou_14_16, in_15_17, ou_15_17 );
  u   u_15_18( clock,enable,reset,set,in_14_18, ou_14_17, in_15_18, ou_15_18 );
  u   u_15_19( clock,enable,reset,set,in_14_19, ou_14_18, in_15_19, ou_15_19 );
  u   u_15_20( clock,enable,reset,set,in_14_20, ou_14_19, in_15_20, ou_15_20 );
  u   u_15_21( clock,enable,reset,set,in_14_21, ou_14_20, in_15_21, ou_15_21 );
  u   u_15_22( clock,enable,reset,set,in_14_22, ou_14_21, in_15_22, ou_15_22 );
  u   u_15_23( clock,enable,reset,set,in_14_23, ou_14_22, in_15_23, ou_15_23 );
  u   u_15_24( clock,enable,reset,set,in_14_24, ou_14_23, in_15_24, ou_15_24 );
  u   u_15_25( clock,enable,reset,set,in_14_25, ou_14_24, in_15_25, ou_15_25 );
  u   u_16_01( clock,enable,reset,set,in_15_01, ou_15_00, in_16_01, ou_16_01 );
  u   u_16_02( clock,enable,reset,set,in_15_02, ou_15_01, in_16_02, ou_16_02 );
  u   u_16_03( clock,enable,reset,set,in_15_03, ou_15_02, in_16_03, ou_16_03 );
  u   u_16_04( clock,enable,reset,set,in_15_04, ou_15_03, in_16_04, ou_16_04 );
  u   u_16_05( clock,enable,reset,set,in_15_05, ou_15_04, in_16_05, ou_16_05 );
  u   u_16_06( clock,enable,reset,set,in_15_06, ou_15_05, in_16_06, ou_16_06 );
  u   u_16_07( clock,enable,reset,set,in_15_07, ou_15_06, in_16_07, ou_16_07 );
  u   u_16_08( clock,enable,reset,set,in_15_08, ou_15_07, in_16_08, ou_16_08 );
  u   u_16_09( clock,enable,reset,set,in_15_09, ou_15_08, in_16_09, ou_16_09 );
  u   u_16_10( clock,enable,reset,set,in_15_10, ou_15_09, in_16_10, ou_16_10 );
  u   u_16_11( clock,enable,reset,set,in_15_11, ou_15_10, in_16_11, ou_16_11 );
  u   u_16_12( clock,enable,reset,set,in_15_12, ou_15_11, in_16_12, ou_16_12 );
  u   u_16_13( clock,enable,reset,set,in_15_13, ou_15_12, in_16_13, ou_16_13 );
  u   u_16_14( clock,enable,reset,set,in_15_14, ou_15_13, in_16_14, ou_16_14 );
  u   u_16_15( clock,enable,reset,set,in_15_15, ou_15_14, in_16_15, ou_16_15 );
  u   u_16_16( clock,enable,reset,set,in_15_16, ou_15_15, in_16_16, ou_16_16 );
  u   u_16_17( clock,enable,reset,set,in_15_17, ou_15_16, in_16_17, ou_16_17 );
  u   u_16_18( clock,enable,reset,set,in_15_18, ou_15_17, in_16_18, ou_16_18 );
  u   u_16_19( clock,enable,reset,set,in_15_19, ou_15_18, in_16_19, ou_16_19 );
  u   u_16_20( clock,enable,reset,set,in_15_20, ou_15_19, in_16_20, ou_16_20 );
  u   u_16_21( clock,enable,reset,set,in_15_21, ou_15_20, in_16_21, ou_16_21 );
  u   u_16_22( clock,enable,reset,set,in_15_22, ou_15_21, in_16_22, ou_16_22 );
  u   u_16_23( clock,enable,reset,set,in_15_23, ou_15_22, in_16_23, ou_16_23 );
  u   u_16_24( clock,enable,reset,set,in_15_24, ou_15_23, in_16_24, ou_16_24 );
  u   u_16_25( clock,enable,reset,set,in_15_25, ou_15_24, in_16_25, ou_16_25 );
  u   u_17_01( clock,enable,reset,set,in_16_01, ou_16_00, in_17_01, ou_17_01 );
  u   u_17_02( clock,enable,reset,set,in_16_02, ou_16_01, in_17_02, ou_17_02 );
  u   u_17_03( clock,enable,reset,set,in_16_03, ou_16_02, in_17_03, ou_17_03 );
  u   u_17_04( clock,enable,reset,set,in_16_04, ou_16_03, in_17_04, ou_17_04 );
  u   u_17_05( clock,enable,reset,set,in_16_05, ou_16_04, in_17_05, ou_17_05 );
  u   u_17_06( clock,enable,reset,set,in_16_06, ou_16_05, in_17_06, ou_17_06 );
  u   u_17_07( clock,enable,reset,set,in_16_07, ou_16_06, in_17_07, ou_17_07 );
  u   u_17_08( clock,enable,reset,set,in_16_08, ou_16_07, in_17_08, ou_17_08 );
  u   u_17_09( clock,enable,reset,set,in_16_09, ou_16_08, in_17_09, ou_17_09 );
  u   u_17_10( clock,enable,reset,set,in_16_10, ou_16_09, in_17_10, ou_17_10 );
  u   u_17_11( clock,enable,reset,set,in_16_11, ou_16_10, in_17_11, ou_17_11 );
  u   u_17_12( clock,enable,reset,set,in_16_12, ou_16_11, in_17_12, ou_17_12 );
  u   u_17_13( clock,enable,reset,set,in_16_13, ou_16_12, in_17_13, ou_17_13 );
  u   u_17_14( clock,enable,reset,set,in_16_14, ou_16_13, in_17_14, ou_17_14 );
  u   u_17_15( clock,enable,reset,set,in_16_15, ou_16_14, in_17_15, ou_17_15 );
  u   u_17_16( clock,enable,reset,set,in_16_16, ou_16_15, in_17_16, ou_17_16 );
  u   u_17_17( clock,enable,reset,set,in_16_17, ou_16_16, in_17_17, ou_17_17 );
  u   u_17_18( clock,enable,reset,set,in_16_18, ou_16_17, in_17_18, ou_17_18 );
  u   u_17_19( clock,enable,reset,set,in_16_19, ou_16_18, in_17_19, ou_17_19 );
  u   u_17_20( clock,enable,reset,set,in_16_20, ou_16_19, in_17_20, ou_17_20 );
  u   u_17_21( clock,enable,reset,set,in_16_21, ou_16_20, in_17_21, ou_17_21 );
  u   u_17_22( clock,enable,reset,set,in_16_22, ou_16_21, in_17_22, ou_17_22 );
  u   u_17_23( clock,enable,reset,set,in_16_23, ou_16_22, in_17_23, ou_17_23 );
  u   u_17_24( clock,enable,reset,set,in_16_24, ou_16_23, in_17_24, ou_17_24 );
  u   u_17_25( clock,enable,reset,set,in_16_25, ou_16_24, in_17_25, ou_17_25 );
  u   u_18_01( clock,enable,reset,set,in_17_01, ou_17_00, in_18_01, ou_18_01 );
  u   u_18_02( clock,enable,reset,set,in_17_02, ou_17_01, in_18_02, ou_18_02 );
  u   u_18_03( clock,enable,reset,set,in_17_03, ou_17_02, in_18_03, ou_18_03 );
  u   u_18_04( clock,enable,reset,set,in_17_04, ou_17_03, in_18_04, ou_18_04 );
  u   u_18_05( clock,enable,reset,set,in_17_05, ou_17_04, in_18_05, ou_18_05 );
  u   u_18_06( clock,enable,reset,set,in_17_06, ou_17_05, in_18_06, ou_18_06 );
  u   u_18_07( clock,enable,reset,set,in_17_07, ou_17_06, in_18_07, ou_18_07 );
  u   u_18_08( clock,enable,reset,set,in_17_08, ou_17_07, in_18_08, ou_18_08 );
  u   u_18_09( clock,enable,reset,set,in_17_09, ou_17_08, in_18_09, ou_18_09 );
  u   u_18_10( clock,enable,reset,set,in_17_10, ou_17_09, in_18_10, ou_18_10 );
  u   u_18_11( clock,enable,reset,set,in_17_11, ou_17_10, in_18_11, ou_18_11 );
  u   u_18_12( clock,enable,reset,set,in_17_12, ou_17_11, in_18_12, ou_18_12 );
  u   u_18_13( clock,enable,reset,set,in_17_13, ou_17_12, in_18_13, ou_18_13 );
  u   u_18_14( clock,enable,reset,set,in_17_14, ou_17_13, in_18_14, ou_18_14 );
  u   u_18_15( clock,enable,reset,set,in_17_15, ou_17_14, in_18_15, ou_18_15 );
  u   u_18_16( clock,enable,reset,set,in_17_16, ou_17_15, in_18_16, ou_18_16 );
  u   u_18_17( clock,enable,reset,set,in_17_17, ou_17_16, in_18_17, ou_18_17 );
  u   u_18_18( clock,enable,reset,set,in_17_18, ou_17_17, in_18_18, ou_18_18 );
  u   u_18_19( clock,enable,reset,set,in_17_19, ou_17_18, in_18_19, ou_18_19 );
  u   u_18_20( clock,enable,reset,set,in_17_20, ou_17_19, in_18_20, ou_18_20 );
  u   u_18_21( clock,enable,reset,set,in_17_21, ou_17_20, in_18_21, ou_18_21 );
  u   u_18_22( clock,enable,reset,set,in_17_22, ou_17_21, in_18_22, ou_18_22 );
  u   u_18_23( clock,enable,reset,set,in_17_23, ou_17_22, in_18_23, ou_18_23 );
  u   u_18_24( clock,enable,reset,set,in_17_24, ou_17_23, in_18_24, ou_18_24 );
  u   u_18_25( clock,enable,reset,set,in_17_25, ou_17_24, in_18_25, ou_18_25 );
  u   u_19_01( clock,enable,reset,set,in_18_01, ou_18_00, in_19_01, ou_19_01 );
  u   u_19_02( clock,enable,reset,set,in_18_02, ou_18_01, in_19_02, ou_19_02 );
  u   u_19_03( clock,enable,reset,set,in_18_03, ou_18_02, in_19_03, ou_19_03 );
  u   u_19_04( clock,enable,reset,set,in_18_04, ou_18_03, in_19_04, ou_19_04 );
  u   u_19_05( clock,enable,reset,set,in_18_05, ou_18_04, in_19_05, ou_19_05 );
  u   u_19_06( clock,enable,reset,set,in_18_06, ou_18_05, in_19_06, ou_19_06 );
  u   u_19_07( clock,enable,reset,set,in_18_07, ou_18_06, in_19_07, ou_19_07 );
  u   u_19_08( clock,enable,reset,set,in_18_08, ou_18_07, in_19_08, ou_19_08 );
  u   u_19_09( clock,enable,reset,set,in_18_09, ou_18_08, in_19_09, ou_19_09 );
  u   u_19_10( clock,enable,reset,set,in_18_10, ou_18_09, in_19_10, ou_19_10 );
  u   u_19_11( clock,enable,reset,set,in_18_11, ou_18_10, in_19_11, ou_19_11 );
  u   u_19_12( clock,enable,reset,set,in_18_12, ou_18_11, in_19_12, ou_19_12 );
  u   u_19_13( clock,enable,reset,set,in_18_13, ou_18_12, in_19_13, ou_19_13 );
  u   u_19_14( clock,enable,reset,set,in_18_14, ou_18_13, in_19_14, ou_19_14 );
  u   u_19_15( clock,enable,reset,set,in_18_15, ou_18_14, in_19_15, ou_19_15 );
  u   u_19_16( clock,enable,reset,set,in_18_16, ou_18_15, in_19_16, ou_19_16 );
  u   u_19_17( clock,enable,reset,set,in_18_17, ou_18_16, in_19_17, ou_19_17 );
  u   u_19_18( clock,enable,reset,set,in_18_18, ou_18_17, in_19_18, ou_19_18 );
  u   u_19_19( clock,enable,reset,set,in_18_19, ou_18_18, in_19_19, ou_19_19 );
  u   u_19_20( clock,enable,reset,set,in_18_20, ou_18_19, in_19_20, ou_19_20 );
  u   u_19_21( clock,enable,reset,set,in_18_21, ou_18_20, in_19_21, ou_19_21 );
  u   u_19_22( clock,enable,reset,set,in_18_22, ou_18_21, in_19_22, ou_19_22 );
  u   u_19_23( clock,enable,reset,set,in_18_23, ou_18_22, in_19_23, ou_19_23 );
  u   u_19_24( clock,enable,reset,set,in_18_24, ou_18_23, in_19_24, ou_19_24 );
  u   u_19_25( clock,enable,reset,set,in_18_25, ou_18_24, in_19_25, ou_19_25 );
  u   u_20_01( clock,enable,reset,set,in_19_01, ou_19_00, in_20_01, ou_20_01 );
  u   u_20_02( clock,enable,reset,set,in_19_02, ou_19_01, in_20_02, ou_20_02 );
  u   u_20_03( clock,enable,reset,set,in_19_03, ou_19_02, in_20_03, ou_20_03 );
  u   u_20_04( clock,enable,reset,set,in_19_04, ou_19_03, in_20_04, ou_20_04 );
  u   u_20_05( clock,enable,reset,set,in_19_05, ou_19_04, in_20_05, ou_20_05 );
  u   u_20_06( clock,enable,reset,set,in_19_06, ou_19_05, in_20_06, ou_20_06 );
  u   u_20_07( clock,enable,reset,set,in_19_07, ou_19_06, in_20_07, ou_20_07 );
  u   u_20_08( clock,enable,reset,set,in_19_08, ou_19_07, in_20_08, ou_20_08 );
  u   u_20_09( clock,enable,reset,set,in_19_09, ou_19_08, in_20_09, ou_20_09 );
  u   u_20_10( clock,enable,reset,set,in_19_10, ou_19_09, in_20_10, ou_20_10 );
  u   u_20_11( clock,enable,reset,set,in_19_11, ou_19_10, in_20_11, ou_20_11 );
  u   u_20_12( clock,enable,reset,set,in_19_12, ou_19_11, in_20_12, ou_20_12 );
  u   u_20_13( clock,enable,reset,set,in_19_13, ou_19_12, in_20_13, ou_20_13 );
  u   u_20_14( clock,enable,reset,set,in_19_14, ou_19_13, in_20_14, ou_20_14 );
  u   u_20_15( clock,enable,reset,set,in_19_15, ou_19_14, in_20_15, ou_20_15 );
  u   u_20_16( clock,enable,reset,set,in_19_16, ou_19_15, in_20_16, ou_20_16 );
  u   u_20_17( clock,enable,reset,set,in_19_17, ou_19_16, in_20_17, ou_20_17 );
  u   u_20_18( clock,enable,reset,set,in_19_18, ou_19_17, in_20_18, ou_20_18 );
  u   u_20_19( clock,enable,reset,set,in_19_19, ou_19_18, in_20_19, ou_20_19 );
  u   u_20_20( clock,enable,reset,set,in_19_20, ou_19_19, in_20_20, ou_20_20 );
  u   u_20_21( clock,enable,reset,set,in_19_21, ou_19_20, in_20_21, ou_20_21 );
  u   u_20_22( clock,enable,reset,set,in_19_22, ou_19_21, in_20_22, ou_20_22 );
  u   u_20_23( clock,enable,reset,set,in_19_23, ou_19_22, in_20_23, ou_20_23 );
  u   u_20_24( clock,enable,reset,set,in_19_24, ou_19_23, in_20_24, ou_20_24 );
  u   u_20_25( clock,enable,reset,set,in_19_25, ou_19_24, in_20_25, ou_20_25 );
  u   u_21_01( clock,enable,reset,set,in_20_01, ou_20_00, in_21_01, ou_21_01 );
  u   u_21_02( clock,enable,reset,set,in_20_02, ou_20_01, in_21_02, ou_21_02 );
  u   u_21_03( clock,enable,reset,set,in_20_03, ou_20_02, in_21_03, ou_21_03 );
  u   u_21_04( clock,enable,reset,set,in_20_04, ou_20_03, in_21_04, ou_21_04 );
  u   u_21_05( clock,enable,reset,set,in_20_05, ou_20_04, in_21_05, ou_21_05 );
  u   u_21_06( clock,enable,reset,set,in_20_06, ou_20_05, in_21_06, ou_21_06 );
  u   u_21_07( clock,enable,reset,set,in_20_07, ou_20_06, in_21_07, ou_21_07 );
  u   u_21_08( clock,enable,reset,set,in_20_08, ou_20_07, in_21_08, ou_21_08 );
  u   u_21_09( clock,enable,reset,set,in_20_09, ou_20_08, in_21_09, ou_21_09 );
  u   u_21_10( clock,enable,reset,set,in_20_10, ou_20_09, in_21_10, ou_21_10 );
  u   u_21_11( clock,enable,reset,set,in_20_11, ou_20_10, in_21_11, ou_21_11 );
  u   u_21_12( clock,enable,reset,set,in_20_12, ou_20_11, in_21_12, ou_21_12 );
  u   u_21_13( clock,enable,reset,set,in_20_13, ou_20_12, in_21_13, ou_21_13 );
  u   u_21_14( clock,enable,reset,set,in_20_14, ou_20_13, in_21_14, ou_21_14 );
  u   u_21_15( clock,enable,reset,set,in_20_15, ou_20_14, in_21_15, ou_21_15 );
  u   u_21_16( clock,enable,reset,set,in_20_16, ou_20_15, in_21_16, ou_21_16 );
  u   u_21_17( clock,enable,reset,set,in_20_17, ou_20_16, in_21_17, ou_21_17 );
  u   u_21_18( clock,enable,reset,set,in_20_18, ou_20_17, in_21_18, ou_21_18 );
  u   u_21_19( clock,enable,reset,set,in_20_19, ou_20_18, in_21_19, ou_21_19 );
  u   u_21_20( clock,enable,reset,set,in_20_20, ou_20_19, in_21_20, ou_21_20 );
  u   u_21_21( clock,enable,reset,set,in_20_21, ou_20_20, in_21_21, ou_21_21 );
  u   u_21_22( clock,enable,reset,set,in_20_22, ou_20_21, in_21_22, ou_21_22 );
  u   u_21_23( clock,enable,reset,set,in_20_23, ou_20_22, in_21_23, ou_21_23 );
  u   u_21_24( clock,enable,reset,set,in_20_24, ou_20_23, in_21_24, ou_21_24 );
  u   u_21_25( clock,enable,reset,set,in_20_25, ou_20_24, in_21_25, ou_21_25 );
  u   u_22_01( clock,enable,reset,set,in_21_01, ou_21_00, in_22_01, ou_22_01 );
  u   u_22_02( clock,enable,reset,set,in_21_02, ou_21_01, in_22_02, ou_22_02 );
  u   u_22_03( clock,enable,reset,set,in_21_03, ou_21_02, in_22_03, ou_22_03 );
  u   u_22_04( clock,enable,reset,set,in_21_04, ou_21_03, in_22_04, ou_22_04 );
  u   u_22_05( clock,enable,reset,set,in_21_05, ou_21_04, in_22_05, ou_22_05 );
  u   u_22_06( clock,enable,reset,set,in_21_06, ou_21_05, in_22_06, ou_22_06 );
  u   u_22_07( clock,enable,reset,set,in_21_07, ou_21_06, in_22_07, ou_22_07 );
  u   u_22_08( clock,enable,reset,set,in_21_08, ou_21_07, in_22_08, ou_22_08 );
  u   u_22_09( clock,enable,reset,set,in_21_09, ou_21_08, in_22_09, ou_22_09 );
  u   u_22_10( clock,enable,reset,set,in_21_10, ou_21_09, in_22_10, ou_22_10 );
  u   u_22_11( clock,enable,reset,set,in_21_11, ou_21_10, in_22_11, ou_22_11 );
  u   u_22_12( clock,enable,reset,set,in_21_12, ou_21_11, in_22_12, ou_22_12 );
  u   u_22_13( clock,enable,reset,set,in_21_13, ou_21_12, in_22_13, ou_22_13 );
  u   u_22_14( clock,enable,reset,set,in_21_14, ou_21_13, in_22_14, ou_22_14 );
  u   u_22_15( clock,enable,reset,set,in_21_15, ou_21_14, in_22_15, ou_22_15 );
  u   u_22_16( clock,enable,reset,set,in_21_16, ou_21_15, in_22_16, ou_22_16 );
  u   u_22_17( clock,enable,reset,set,in_21_17, ou_21_16, in_22_17, ou_22_17 );
  u   u_22_18( clock,enable,reset,set,in_21_18, ou_21_17, in_22_18, ou_22_18 );
  u   u_22_19( clock,enable,reset,set,in_21_19, ou_21_18, in_22_19, ou_22_19 );
  u   u_22_20( clock,enable,reset,set,in_21_20, ou_21_19, in_22_20, ou_22_20 );
  u   u_22_21( clock,enable,reset,set,in_21_21, ou_21_20, in_22_21, ou_22_21 );
  u   u_22_22( clock,enable,reset,set,in_21_22, ou_21_21, in_22_22, ou_22_22 );
  u   u_22_23( clock,enable,reset,set,in_21_23, ou_21_22, in_22_23, ou_22_23 );
  u   u_22_24( clock,enable,reset,set,in_21_24, ou_21_23, in_22_24, ou_22_24 );
  u   u_22_25( clock,enable,reset,set,in_21_25, ou_21_24, in_22_25, ou_22_25 );
  u   u_23_01( clock,enable,reset,set,in_22_01, ou_22_00, in_23_01, ou_23_01 );
  u   u_23_02( clock,enable,reset,set,in_22_02, ou_22_01, in_23_02, ou_23_02 );
  u   u_23_03( clock,enable,reset,set,in_22_03, ou_22_02, in_23_03, ou_23_03 );
  u   u_23_04( clock,enable,reset,set,in_22_04, ou_22_03, in_23_04, ou_23_04 );
  u   u_23_05( clock,enable,reset,set,in_22_05, ou_22_04, in_23_05, ou_23_05 );
  u   u_23_06( clock,enable,reset,set,in_22_06, ou_22_05, in_23_06, ou_23_06 );
  u   u_23_07( clock,enable,reset,set,in_22_07, ou_22_06, in_23_07, ou_23_07 );
  u   u_23_08( clock,enable,reset,set,in_22_08, ou_22_07, in_23_08, ou_23_08 );
  u   u_23_09( clock,enable,reset,set,in_22_09, ou_22_08, in_23_09, ou_23_09 );
  u   u_23_10( clock,enable,reset,set,in_22_10, ou_22_09, in_23_10, ou_23_10 );
  u   u_23_11( clock,enable,reset,set,in_22_11, ou_22_10, in_23_11, ou_23_11 );
  u   u_23_12( clock,enable,reset,set,in_22_12, ou_22_11, in_23_12, ou_23_12 );
  u   u_23_13( clock,enable,reset,set,in_22_13, ou_22_12, in_23_13, ou_23_13 );
  u   u_23_14( clock,enable,reset,set,in_22_14, ou_22_13, in_23_14, ou_23_14 );
  u   u_23_15( clock,enable,reset,set,in_22_15, ou_22_14, in_23_15, ou_23_15 );
  u   u_23_16( clock,enable,reset,set,in_22_16, ou_22_15, in_23_16, ou_23_16 );
  u   u_23_17( clock,enable,reset,set,in_22_17, ou_22_16, in_23_17, ou_23_17 );
  u   u_23_18( clock,enable,reset,set,in_22_18, ou_22_17, in_23_18, ou_23_18 );
  u   u_23_19( clock,enable,reset,set,in_22_19, ou_22_18, in_23_19, ou_23_19 );
  u   u_23_20( clock,enable,reset,set,in_22_20, ou_22_19, in_23_20, ou_23_20 );
  u   u_23_21( clock,enable,reset,set,in_22_21, ou_22_20, in_23_21, ou_23_21 );
  u   u_23_22( clock,enable,reset,set,in_22_22, ou_22_21, in_23_22, ou_23_22 );
  u   u_23_23( clock,enable,reset,set,in_22_23, ou_22_22, in_23_23, ou_23_23 );
  u   u_23_24( clock,enable,reset,set,in_22_24, ou_22_23, in_23_24, ou_23_24 );
  u   u_23_25( clock,enable,reset,set,in_22_25, ou_22_24, in_23_25, ou_23_25 );
  u   u_24_01( clock,enable,reset,set,in_23_01, ou_23_00, in_24_01, ou_24_01 );
  u   u_24_02( clock,enable,reset,set,in_23_02, ou_23_01, in_24_02, ou_24_02 );
  u   u_24_03( clock,enable,reset,set,in_23_03, ou_23_02, in_24_03, ou_24_03 );
  u   u_24_04( clock,enable,reset,set,in_23_04, ou_23_03, in_24_04, ou_24_04 );
  u   u_24_05( clock,enable,reset,set,in_23_05, ou_23_04, in_24_05, ou_24_05 );
  u   u_24_06( clock,enable,reset,set,in_23_06, ou_23_05, in_24_06, ou_24_06 );
  u   u_24_07( clock,enable,reset,set,in_23_07, ou_23_06, in_24_07, ou_24_07 );
  u   u_24_08( clock,enable,reset,set,in_23_08, ou_23_07, in_24_08, ou_24_08 );
  u   u_24_09( clock,enable,reset,set,in_23_09, ou_23_08, in_24_09, ou_24_09 );
  u   u_24_10( clock,enable,reset,set,in_23_10, ou_23_09, in_24_10, ou_24_10 );
  u   u_24_11( clock,enable,reset,set,in_23_11, ou_23_10, in_24_11, ou_24_11 );
  u   u_24_12( clock,enable,reset,set,in_23_12, ou_23_11, in_24_12, ou_24_12 );
  u   u_24_13( clock,enable,reset,set,in_23_13, ou_23_12, in_24_13, ou_24_13 );
  u   u_24_14( clock,enable,reset,set,in_23_14, ou_23_13, in_24_14, ou_24_14 );
  u   u_24_15( clock,enable,reset,set,in_23_15, ou_23_14, in_24_15, ou_24_15 );
  u   u_24_16( clock,enable,reset,set,in_23_16, ou_23_15, in_24_16, ou_24_16 );
  u   u_24_17( clock,enable,reset,set,in_23_17, ou_23_16, in_24_17, ou_24_17 );
  u   u_24_18( clock,enable,reset,set,in_23_18, ou_23_17, in_24_18, ou_24_18 );
  u   u_24_19( clock,enable,reset,set,in_23_19, ou_23_18, in_24_19, ou_24_19 );
  u   u_24_20( clock,enable,reset,set,in_23_20, ou_23_19, in_24_20, ou_24_20 );
  u   u_24_21( clock,enable,reset,set,in_23_21, ou_23_20, in_24_21, ou_24_21 );
  u   u_24_22( clock,enable,reset,set,in_23_22, ou_23_21, in_24_22, ou_24_22 );
  u   u_24_23( clock,enable,reset,set,in_23_23, ou_23_22, in_24_23, ou_24_23 );
  u   u_24_24( clock,enable,reset,set,in_23_24, ou_23_23, in_24_24, ou_24_24 );
  u   u_24_25( clock,enable,reset,set,in_23_25, ou_23_24, in_24_25, ou_24_25 );
  u   u_25_01( clock,enable,reset,set,in_24_01, ou_24_00, in_25_01, ou_25_01 );
  u   u_25_02( clock,enable,reset,set,in_24_02, ou_24_01, in_25_02, ou_25_02 );
  u   u_25_03( clock,enable,reset,set,in_24_03, ou_24_02, in_25_03, ou_25_03 );
  u   u_25_04( clock,enable,reset,set,in_24_04, ou_24_03, in_25_04, ou_25_04 );
  u   u_25_05( clock,enable,reset,set,in_24_05, ou_24_04, in_25_05, ou_25_05 );
  u   u_25_06( clock,enable,reset,set,in_24_06, ou_24_05, in_25_06, ou_25_06 );
  u   u_25_07( clock,enable,reset,set,in_24_07, ou_24_06, in_25_07, ou_25_07 );
  u   u_25_08( clock,enable,reset,set,in_24_08, ou_24_07, in_25_08, ou_25_08 );
  u   u_25_09( clock,enable,reset,set,in_24_09, ou_24_08, in_25_09, ou_25_09 );
  u   u_25_10( clock,enable,reset,set,in_24_10, ou_24_09, in_25_10, ou_25_10 );
  u   u_25_11( clock,enable,reset,set,in_24_11, ou_24_10, in_25_11, ou_25_11 );
  u   u_25_12( clock,enable,reset,set,in_24_12, ou_24_11, in_25_12, ou_25_12 );
  u   u_25_13( clock,enable,reset,set,in_24_13, ou_24_12, in_25_13, ou_25_13 );
  u   u_25_14( clock,enable,reset,set,in_24_14, ou_24_13, in_25_14, ou_25_14 );
  u   u_25_15( clock,enable,reset,set,in_24_15, ou_24_14, in_25_15, ou_25_15 );
  u   u_25_16( clock,enable,reset,set,in_24_16, ou_24_15, in_25_16, ou_25_16 );
  u   u_25_17( clock,enable,reset,set,in_24_17, ou_24_16, in_25_17, ou_25_17 );
  u   u_25_18( clock,enable,reset,set,in_24_18, ou_24_17, in_25_18, ou_25_18 );
  u   u_25_19( clock,enable,reset,set,in_24_19, ou_24_18, in_25_19, ou_25_19 );
  u   u_25_20( clock,enable,reset,set,in_24_20, ou_24_19, in_25_20, ou_25_20 );
  u   u_25_21( clock,enable,reset,set,in_24_21, ou_24_20, in_25_21, ou_25_21 );
  u   u_25_22( clock,enable,reset,set,in_24_22, ou_24_21, in_25_22, ou_25_22 );
  u   u_25_23( clock,enable,reset,set,in_24_23, ou_24_22, in_25_23, ou_25_23 );
  u   u_25_24( clock,enable,reset,set,in_24_24, ou_24_23, in_25_24, ou_25_24 );
  u   u_25_25( clock,enable,reset,set,in_24_25, ou_24_24, in_25_25, ou_25_25 );

endmodule
